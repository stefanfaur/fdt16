module ControlUnit(
    input clk, reset,
    input [5:0] opcode,
    input [3:0] flags,
    output reg [4:0] state
);


endmodule